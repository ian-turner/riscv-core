module controlunit(
	// inputs
	input logic [6:0] opcode,
	input logic [2:0] funct3,
	input logic [6:0] funct7,
	input logic [11:0] csr,

	// outputs
	// ...
);

endmodule
