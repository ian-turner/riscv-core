/* Copyright 2020 Jason Bakos, Philip Conrad, Charles Daniels */

/* Top-level module for CSCE611 RISC-V CPU, for running under simulation.  In
 * this case, the I/Os and clock are driven by the simulator. */

module simtop;

	logic clk;
	logic [6:0] HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7;
	logic [3:0] KEY;
	logic [17:0] SW;

	top dut
	(
		//////////// CLOCK //////////
		.CLOCK_50(clk),
		.CLOCK2_50(),
	    	.CLOCK3_50(),

		//////////// LED //////////
		.LEDG(),
		.LEDR(),

		//////////// KEY //////////
		.KEY(KEY),

		//////////// SW //////////
		.SW(SW),

		//////////// SEG7 //////////
		.HEX0(HEX0),
		.HEX1(HEX1),
		.HEX2(HEX2),
		.HEX3(HEX3),
		.HEX4(HEX4),
		.HEX5(HEX5),
		.HEX6(HEX6),
		.HEX7(HEX7)
	);

	logic [31:0] io0_out;
	logic [31:0] io0_in;

	cpu _cpu(clk, KEY[0], io0_in, io0_out);

	// pulse reset (active low)
	initial begin
		KEY <= 4'he;
		#10;
		KEY <= 4'hf;

		// 10 ticks = 1 clock tick

		#1000; // <- 100 clock ticks

		// verify register file
		// we can ignore 0 register because 0 is hard coded in regfile
		for (int i=0; i<32; i++) begin
			$display("register %d: 0x%h", i, _cpu._regfile.mem[i]);
		end
	end
	
	// drive clock
	always begin
		clk <= 1'b0; #5;
		clk <= 1'b1; #5;
	end

	always_comb begin
		io0_in = {14'b0, SW};
	end
	
	// assign simulated switch values
	assign SW = 18'd12345;

endmodule

